module TubeTest

(
	
	input clk,
	input reg Key[3:0],
	input reg Sw[7:0],
	
	output reg Dot,
	output reg Seg[6:0],
	output reg Led[0:7],
	
);

	

	// Module Item(s)

endmodule
